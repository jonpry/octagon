----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:47:22 04/23/2013 
-- Design Name: 
-- Module Name:    octagon - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

use work.octagon_types.all;

entity octagon is
	Port ( 
		clk : in  std_logic;
		jump_target 	: in std_logic_vector(IM_BITS-1 downto 0);
		running 			: in std_logic_vector(7 downto 0);
		int 				: in std_logic_vector(7 downto 0);
		do_jump				: in std_logic;
		notrim_o : out std_logic_vector(20 downto 0);
		routq		: out rfetchout_type;
		alu2outq : out alu2out_type;
		tagidx			: in std_logic_vector(2 downto 0);
		tagadr			: in std_logic_vector(3 downto 0);
		tagval			: in std_logic_vector(IM_BITS-1 downto 10);
		tagwe				: in std_logic;
		imemidx			: in std_logic_vector(2 downto 0);
		imemadr			: in std_logic_vector(7 downto 0);
		imemval			: in std_logic_vector(31 downto 0);
		ipresent			: in std_logic;
		imemwe			: in std_logic;
		reg_we			: in std_logic
	);
end octagon;

architecture Behavioral of octagon is

signal pcin : pcin_type;
signal pcout : pcout_type;
signal icin : icfetchin_type;
signal icout : icfetchout_type;
signal muxout : icmuxout_type;
signal decout : decout_type;
signal rin : rfetchin_type;
signal rout : rfetchout_type;
signal alu1out : alu1out_type;
signal alu2out : alu2out_type;
signal jumpout : jumpout_type;

begin

routq <= rout;
alu2outq <= alu2out;

--1 PC
--2 Tag
--3 Mux
--4 decode
--5 R fetch
--6 alu
--7 alu
--8 alu - jump - load stall - or stall if store still pending
--9 alu
--11 store

pcin.jump_target <= jump_target;
pcin.running <= running;
pcin.int <= int;
pcin.jump <= do_jump;
pcin.valid <= jumpout.valid;

icin.pcout <= pcout;
icin.tagval <= tagval;
icin.tagadr <= tagadr;
icin.tagidx <= tagidx;
icin.tagwe <= tagwe;
icin.imemval <= imemval;
icin.imemadr <= imemadr;
icin.imemidx <= imemidx;
icin.imemwe <= imemwe;
icin.ipresent <= ipresent;

rin.decout <= decout;
rin.reg_val <= imemval;
rin.reg_adr <= imemadr;
rin.reg_we <= reg_we;

pc_module: entity work.pc_module port map(clk,pcin,pcout);  --1
ic_fetch : entity work.ic_fetch port map(clk,icin,icout);	--2
ic_mux : entity work.ic_mux port map(clk,icout,muxout);		--3
decode : entity work.decode port map(clk,muxout,decout);		--4
r_fetch : entity work.r_fetch port map(clk,rin,rout);			--5
alu1 : entity work.alu1 port map(clk,rout,alu1out);			--6
alu2 : entity work.alu2 port map(clk,alu1out,alu2out);		--7
jump : entity work.jump port map(clk,alu2out,jumpout);		--8

process(clk)
variable notrim : std_logic_vector(20 downto 0);
begin
	if clk='1' and clk'Event then
		notrim := (others => '0');
		notrim(4 downto 0) := notrim(4 downto 0) or decout.r_dest;
		notrim(11 downto 10) := notrim(11 downto 10) or decout.memsize;
		notrim(15) := notrim(15) or decout.link;
		notrim(16) := notrim(16) or decout.rfe;
		notrim(16) := notrim(16) or decout.load;
		notrim(17) := notrim(17) or decout.store;
		notrim(17) := notrim(17) or decout.load_unsigned;
		notrim(18) := notrim(18) or decout.arith;
		notrim(18) := notrim(18) or decout.slt;
		notrim(19) := notrim(19) or decout.logic;
		notrim(20) := notrim(20) or decout.jump;
		notrim(20) := notrim(20) or decout.math_unsigned;

		notrim_o <= notrim;


	end if;
end process;

end Behavioral;

